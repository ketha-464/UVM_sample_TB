//interface
interface our_interface(input logic clk);

  //input_1;
  //input-2;
  logic [7:0]input_1;
  logic [7:0]input_2;
  
  //output_1;
  //output_2;
  logic [15:0]output_1;
  logic [15:0]output_2;
endinterface